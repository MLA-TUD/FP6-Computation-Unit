library ieee;
use ieee.std_logic_1164.all;


entity controller is	
	
end controller;

architecture behavior of controller is
begin	
end behavior;
