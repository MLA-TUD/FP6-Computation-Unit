library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity matrix_multiplier is	
end matrix_multiplier;

architecture behavior of matrix_multiplier is
begin
	
end behavior;
