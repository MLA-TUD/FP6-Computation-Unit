library ieee;
use ieee.std_logic_1164.all;

entity sa_tb is -- systolic array testbench
end sa_tb;

architecture test of sa_tb is
	
	-- ?
begin
	
	process begin
		-- ?
		wait;
	end process;
end test;
