library ieee;
use ieee.std_logic_1164.all;

entity ksa is -- kogge-stone adder
	port ( -- s: sum
		a : in std_logic_vector(7 downto 0);
		b : in std_logic_vector(7 downto 0);
		s : out std_logic_vector(7 downto 0)
	);
end ksa;

architecture behavior of ksa is
	-- ?
begin
	-- ?
end behavior;